library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity circuiteria is
  port(
    clk         : in  std_logic;
    reset       : in  std_logic;
    SDA         : in  std_logic;
    Hab_Dir     : in  std_logic;
    Hab_Dat     : in  std_logic;
    Direccion   : in  std_logic_vector(6 downto 0);
    soy         : out std_logic;
    fin_dato    : out std_logic
  );
end entity circuiteria;

architecture Behavioral of circuiteria is
  signal address_shift_reg : std_logic_vector(6 downto 0) := (others => '0');
  signal data_shift_reg    : std_logic_vector(7 downto 0) := (others => '0');
  signal bit_counter       : integer range 0 to 7 := 0;
begin
  process(clk, reset)
  begin
    if reset = '1' then
      address_shift_reg <= (others => '0');
      data_shift_reg <= (others => '0');
      soy <= '0';
      fin_dato <= '0';
      bit_counter <= 0;
      
    elsif rising_edge(clk) then
      if Hab_Dir = '1' then
        fin_dato <= '0';
        if bit_counter < 7 then
          address_shift_reg <= address_shift_reg(5 downto 0) & SDA;
          bit_counter <= bit_counter + 1;
        else
          if address_shift_reg = Direccion then
            soy <= '1';
          else
            soy <= '0';
          end if;
          bit_counter <= 0;
        end if;

      elsif Hab_Dat = '1' then
        soy <= '0';
        if bit_counter < 8 then
          data_shift_reg <= data_shift_reg(6 downto 0) & SDA;
          bit_counter <= bit_counter + 1;
        else
          fin_dato <= '1';
          bit_counter <= 0;
        end if;

      else
        soy <= '0';
        fin_dato <= '0';
        bit_counter <= 0;
      end if;
    end if;
  end process;
end architecture Behavioral;

