library verilog;
use verilog.vl_types.all;
entity PARTE_A_vlg_check_tst is
    port(
        LED             : in     vl_logic;
        sampler_rx      : in     vl_logic
    );
end PARTE_A_vlg_check_tst;
