library verilog;
use verilog.vl_types.all;
entity PARTE_A_vlg_vec_tst is
end PARTE_A_vlg_vec_tst;
