library verilog;
use verilog.vl_types.all;
entity Circuito_Final_vlg_vec_tst is
end Circuito_Final_vlg_vec_tst;
