library verilog;
use verilog.vl_types.all;
entity PARTE_E_vlg_vec_tst is
end PARTE_E_vlg_vec_tst;
