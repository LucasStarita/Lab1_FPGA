library verilog;
use verilog.vl_types.all;
entity Division_vlg_vec_tst is
end Division_vlg_vec_tst;
