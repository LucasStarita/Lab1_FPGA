library verilog;
use verilog.vl_types.all;
entity PARTE_C_vlg_vec_tst is
end PARTE_C_vlg_vec_tst;
