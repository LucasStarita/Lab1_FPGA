library verilog;
use verilog.vl_types.all;
entity PARTE_C_vlg_check_tst is
    port(
        B               : in     vl_logic;
        C0              : in     vl_logic;
        C1              : in     vl_logic;
        C2              : in     vl_logic;
        C3              : in     vl_logic;
        Z               : in     vl_logic;
        sampler_rx      : in     vl_logic
    );
end PARTE_C_vlg_check_tst;
