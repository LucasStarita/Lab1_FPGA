-- Copyright (C) 1991-2013 Altera Corporation
-- Your use of Altera Corporation's design tools, logic functions 
-- and other software and tools, and its AMPP partner logic 
-- functions, and any output files from any of the foregoing 
-- (including device programming or simulation files), and any 
-- associated documentation or information are expressly subject 
-- to the terms and conditions of the Altera Program License 
-- Subscription Agreement, Altera MegaCore Function License 
-- Agreement, or other applicable license agreement, including, 
-- without limitation, that your use is for the sole purpose of 
-- programming logic devices manufactured by Altera and sold by 
-- Altera or its authorized distributors.  Please refer to the 
-- applicable agreement for further details.

-- Generated by Quartus II Version 13.0.1 Build 232 06/12/2013 Service Pack 1 SJ Web Edition
-- Created on Fri Nov 01 16:02:41 2024

LIBRARY ieee;
USE ieee.std_logic_1164.all;

ENTITY PARTE_E IS
    PORT (
        clock : IN STD_LOGIC;
        reset : IN STD_LOGIC := '0';
        SDA : IN STD_LOGIC := '0';
        fin_dir : IN STD_LOGIC := '0';
        soy : IN STD_LOGIC := '0';
        fin_dato : IN STD_LOGIC := '0';
        Hab_Dir : OUT STD_LOGIC;
        Hab_Dat : OUT STD_LOGIC;
        Hab_ACK : OUT STD_LOGIC
    );
END PARTE_E;

ARCHITECTURE BEHAVIOR OF PARTE_E IS
    TYPE type_fstate IS (Oscioso,Start,Guarda_Direccion,R_W,ACK,Guarda_Dato);
    SIGNAL fstate : type_fstate;
    SIGNAL reg_fstate : type_fstate;
BEGIN
    PROCESS (clock,reg_fstate)
    BEGIN
        IF (clock='1' AND clock'event) THEN
            fstate <= reg_fstate;
        END IF;
    END PROCESS;

    PROCESS (fstate,reset,SDA,fin_dir,soy,fin_dato)
    BEGIN
        IF (reset='1') THEN
            reg_fstate <= Oscioso;
            Hab_Dir <= '0';
            Hab_Dat <= '0';
            Hab_ACK <= '0';
        ELSE
            Hab_Dir <= '0';
            Hab_Dat <= '0';
            Hab_ACK <= '0';
            CASE fstate IS
                WHEN Oscioso =>
                    IF ((SDA = '1')) THEN
                        reg_fstate <= Oscioso;
                    ELSIF ((SDA = '0')) THEN
                        reg_fstate <= Start;
                    -- Inserting 'else' block to prevent latch inference
                    ELSE
                        reg_fstate <= Oscioso;
                    END IF;

                    Hab_ACK <= '0';

                    Hab_Dir <= '0';

                    Hab_Dat <= '0';
                WHEN Start =>
                    reg_fstate <= Guarda_Direccion;

                    Hab_ACK <= '0';

                    Hab_Dir <= '0';

                    Hab_Dat <= '0';
                WHEN Guarda_Direccion =>
                    IF (((fin_dir = '1') AND (soy = '0'))) THEN
                        reg_fstate <= Oscioso;
                    ELSIF (((fin_dir = '1') AND (soy = '1'))) THEN
                        reg_fstate <= R_W;
                    ELSIF ((fin_dir = '0')) THEN
                        reg_fstate <= Guarda_Direccion;
                    -- Inserting 'else' block to prevent latch inference
                    ELSE
                        reg_fstate <= Guarda_Direccion;
                    END IF;

                    Hab_ACK <= '0';

                    Hab_Dir <= '1';

                    Hab_Dat <= '0';
                WHEN R_W =>
                    reg_fstate <= ACK;

                    Hab_ACK <= '0';

                    Hab_Dir <= '0';

                    Hab_Dat <= '0';
                WHEN ACK =>
                    reg_fstate <= Guarda_Dato;

                    Hab_ACK <= '1';

                    Hab_Dir <= '0';

                    Hab_Dat <= '0';
                WHEN Guarda_Dato =>
                    IF ((fin_dato = '0')) THEN
                        reg_fstate <= Guarda_Dato;
                    ELSIF ((fin_dato = '1')) THEN
                        reg_fstate <= Oscioso;
                    -- Inserting 'else' block to prevent latch inference
                    ELSE
                        reg_fstate <= Guarda_Dato;
                    END IF;

                    Hab_ACK <= '0';

                    Hab_Dir <= '0';

                    Hab_Dat <= '1';
                WHEN OTHERS => 
                    Hab_Dir <= 'X';
                    Hab_Dat <= 'X';
                    Hab_ACK <= 'X';
                    report "Reach undefined state";
            END CASE;
        END IF;
    END PROCESS;
END BEHAVIOR;
